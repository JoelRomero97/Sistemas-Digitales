module contadordecada ( 
	e,
	clk,
	clr,
	u,
	d
	) ;

input [1:0] e;
input  clk;
input  clr;
inout [3:0] u;
inout [2:0] d;
