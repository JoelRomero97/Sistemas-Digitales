module marquesina ( 
	e,
	clr,
	clk,
	display,
	sel
	) ;

input [2:0] e;
input  clr;
input  clk;
inout [6:0] display;
inout [2:0] sel;
