module practica6dado ( 
	clear,
	clock,
	enable,
	display
	) ;

input  clear;
input  clock;
input  enable;
inout [6:0] display;
