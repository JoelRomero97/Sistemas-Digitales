module prac52 ( 
	clr,
	clk,
	e,
	l,
	ud,
	d,
	q
	) ;

input  clr;
input  clk;
input  e;
input  l;
input  ud;
input [4:0] d;
inout [4:0] q;
