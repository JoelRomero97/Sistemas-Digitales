module practica6_b_contadorhexadecimal ( 
	clock,
	clear,
	enable,
	display
	) ;

input  clock;
input  clear;
input  enable;
inout [6:0] display;
