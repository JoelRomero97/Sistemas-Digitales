module practica6_d_boleta_contador ( 
	clock,
	clear,
	enable,
	display
	) ;

input  clock;
input  clear;
input  enable;
inout [6:0] display;
