module practica6_c_2_mi_nombre_usando_contador ( 
	clock,
	clear,
	enable,
	display
	) ;

input  clock;
input  clear;
input  enable;
inout [6:0] display;
