module practica5_b_contadorgenerico ( 
	q,
	clock,
	clear,
	enable
	) ;

inout [9:0] q;
input  clock;
input  clear;
input  enable;
