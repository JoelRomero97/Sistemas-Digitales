module practica3 ( 
	x,
	clk,
	clr,
	an0,
	dis
	) ;

input  x;
input  clk;
input  clr;
inout  an0;
inout [6:0] dis;
