LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Sensores IS PORT
(
	CLK, CLR : IN STD_LOGIC;											--CLOCK Y CLEAR
	DISPLAY : OUT STD_LOGIC_VECTOR (6 DOWNTO 0);						--DISPLAY DE 7 SEGMENTOS
	UNI : IN STD_LOGIC_VECTOR (3 DOWNTO 0);								--SALIDA DE CONTADOR DECADA
	DEC : IN STD_LOGIC_VECTOR (2 DOWNTO 0);								--SALIDA DE CONTADOR DECADA
	SEL : STD_LOGIC_VECTOR (2 DOWNTO 0)									--SELECTOR DE MUX
);

ATTRIBUTE PIN_NUMBERS OF Sensores : ENTITY IS
	"DISPLAY(0):21 DISPLAY(1):20 DISPLAY(2):19 DISPLAY(3):18 DISPLAY(4):17 DISPLAY(5):16 DISPLAY(6):15 " &
	"UNI(0):11 UNI(1):10 UNI(2):9 UNI(3):8 " &
	"DEC(0):7 DEC(1):6 DEC(2):5 " &
	"CLR:2 " &
	"SEL(0):14 SEL(1):23 SEL(2):22 ";
END Sensores;

ARCHITECTURE A_Sensores OF Sensores IS
	CONSTANT E1 : STD_LOGIC_VECTOR (3 DOWNTO 0) := '0'&DEC;				--E1 DEL MULTIPLEXOR
	SIGNAL E2 : STD_LOGIC_VECTOR (3 DOWNTO 0) := "0000";				--E2 DEL MULTIPLEXOR
	SIGNAL AN : STD_LOGIC_VECTOR (2 DOWNTO 0);							--ANILLO PARA CONTADOR
	SIGNAL BCD : STD_LOGIC_VECTOR (3 DOWNTO 0);							--SALIDA DE MULTIPLEXOR
BEGIN

		--CONTADOR DE ANILLO
		ContadorAnillo : PROCESS (CLK, CLR)
		BEGIN 
				IF (CLR = '1') THEN
					AN <= "110";
				ELSIF (CLK'EVENT AND CLK = '1') THEN
					CASE AN IS
						WHEN "110" => AN <= "101";
						WHEN "101" => AN <= "011";
						WHEN "011" => AN <= "110";
						WHEN OTHERS => AN <= "---";
					END CASE;
				END IF;
		END PROCESS ContadorAnillo;

		--MULTIPLEXOR
		Multiplexor : PROCESS (BCD, UNI, DEC, E2, AN)
		BEGIN
				SEL <= AN;
				IF (SEL = "110") THEN 
					BCD <= UNI;
				ELSIF (SEL = "101") THEN
					BCD <= E1;
				ELSIF (SEL = "011") THEN
					BCD <= E2;
				ELSE 
					BCD <= "----";
				END IF;
		END PROCESS Multiplexor;

		--CONVERTIDOR DE C�DIGO
		Convertidor : PROCESS (BCD)
		BEGIN
				CASE BCD IS
						WHEN "0000" => DISPLAY <= "0000001";		--0
						WHEN "0001" => DISPLAY <= "1001111";		--1
						WHEN "0010" => DISPLAY <= "0010010";		--2
						WHEN "0011" => DISPLAY <= "0000110";		--3
						WHEN "0100" => DISPLAY <= "1001100";		--4
						WHEN "0101" => DISPLAY <= "0100100";		--5
						WHEN "0110" => DISPLAY <= "0100000";		--6
						WHEN "0111" => DISPLAY <= "0001111";		--7
						WHEN "1000" => DISPLAY <= "0000000";		--8
						WHEN "1001" => DISPLAY <= "0000100";		--9
						WHEN OTHERS => DISPLAY <= "-------";
				END CASE;
		END PROCESS Convertidor; 
END A_Sensores;