module contador ( 
	clr,
	clk,
	e,
	q
	) ;

input  clr;
input  clk;
input  e;
inout [9:0] q;
