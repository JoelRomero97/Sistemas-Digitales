module gal2 ( 
	selector,
	display,
	e0,
	e1,
	clk,
	clr
	) ;

inout [2:0] selector;
inout [6:0] display;
input [3:0] e0;
input [2:0] e1;
input  clk;
input  clr;
