module marquesina ( 
	e,
	clr,
	clk,
	display
	) ;

input [2:0] e;
input  clr;
input  clk;
inout [9:0] display;
