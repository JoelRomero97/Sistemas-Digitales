module sensores ( 
	u,
	d,
	e,
	clr,
	clk
	) ;

inout [3:0] u;
inout [2:0] d;
input [1:0] e;
input  clr;
input  clk;
