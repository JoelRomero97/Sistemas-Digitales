module prac51 ( 
	clr,
	clk,
	e,
	q
	) ;

input  clr;
input  clk;
input  e;
inout [6:0] q;
