module moore ( 
	l,
	clk,
	clr,
	display,
	q,
	teclado
	) ;

input  l;
input  clk;
input  clr;
inout [6:0] display;
inout [2:0] q;
input [3:0] teclado;
