module practica4 ( 
	clr,
	clk,
	display,
	anodo
	) ;

input  clr;
input  clk;
inout [6:0] display;
inout [2:0] anodo;
