module marquesinarom2 ( 
	clr,
	clk,
	dir,
	display,
	an
	) ;

input  clr;
input  clk;
input [3:0] dir;
inout [6:0] display;
inout [2:0] an;
