module prac2 ( 
	clr,
	clk,
	es,
	d,
	q,
	op
	) ;

input  clr;
input  clk;
input  es;
input [6:0] d;
inout [6:0] q;
input [1:0] op;
