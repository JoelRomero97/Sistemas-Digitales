module practica3 ( 
	clear,
	clk,
	x,
	an,
	display
	) ;

input  clear;
input  clk;
input  x;
inout  an;
inout [6:0] display;
