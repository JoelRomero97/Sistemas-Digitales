module marquesinarom1 ( 
	clr,
	clk,
	dir,
	display,
	an
	) ;

input  clr;
input  clk;
input [2:0] dir;
inout [6:0] display;
inout [2:0] an;
