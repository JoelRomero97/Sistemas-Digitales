module practica6_c_mensaje_con_contador ( 
	clock,
	clear,
	enable,
	display
	) ;

input  clock;
input  clear;
input  enable;
inout [6:0] display;
